LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
use ieee.numeric_std.all;
use STD.textio.all;
use ieee.std_logic_textio.all;
use std.env.finish;

 
ENTITY MatrixModulator_tb IS
END MatrixModulator_tb;

architecture Behavioral of MatrixModulator_tb is
    begin
    
end;