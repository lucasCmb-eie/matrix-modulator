library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity MatrixModulator_top is
    port (
        clk   : in std_logic;
        reset : in std_logic );
end entity;

architecture Behavioral of MatrixModulator_top is

begin

    

end architecture;
